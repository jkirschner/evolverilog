module scootBot(output0,output1,output2,output3,input0,input1,input2,input3,input4);

	output output0,output1,output2,output3;
	input input0,input1,input2,input3,input4;
	and #50 (output0_branch0100,input0,input0);
	not #50 (output0_branch0101,input1);
	nand #50 (output0_branch010,output0_branch0100,output0_branch0101);
	and #50 (output0_branch0111010000,input0,input0);
	nand #50 (output0_branch01110100010,input0,input4);
	not #50 (output0_branch011101000110,input1);
	not #50 (output0_branch0111010001110,input1);
	not #50 (output0_branch0111010001111100,input1);
	nand #50 (output0_branch011101000111110,output0_branch0111010001111100,input3);
	and #50 (output0_branch01110100011111,output0_branch011101000111110,input3);
	or #50 (output0_branch0111010001111,input0,output0_branch01110100011111);
	and #50 (output0_branch011101000111,output0_branch0111010001110,output0_branch0111010001111);
	and #50 (output0_branch01110100011,output0_branch011101000110,output0_branch011101000111);
	xor #50 (output0_branch0111010001,output0_branch01110100010,output0_branch01110100011);
	nand #50 (output0_branch011101000,output0_branch0111010000,output0_branch0111010001);
	not #50 (output0_branch011101001101000,input1);
	or #50 (output0_branch011101001101001,input4,input4);
	xor #50 (output0_branch01110100110100,output0_branch011101001101000,output0_branch011101001101001);
	not #50 (output0_branch011101001101010,input0);
	xor #50 (output0_branch01110100110101,output0_branch011101001101010,input3);
	and #50 (output0_branch0111010011010,output0_branch01110100110100,output0_branch01110100110101);
	xor #50 (output0_branch011101001101,output0_branch0111010011010,input0);
	and #50 (output0_branch01110100110,input0,output0_branch011101001101);
	or #50 (output0_branch0111010011,output0_branch01110100110,input0);
	xor #50 (output0_branch011101001,input2,output0_branch0111010011);
	and #50 (output0_branch01110100,output0_branch011101000,output0_branch011101001);
	nand #50 (output0_branch01110101000,input0,input4);
	not #50 (output0_branch011101010010,input1);
	not #50 (output0_branch0111010100110,input1);
	not #50 (output0_branch01110101001111010,input1);
	not #50 (output0_branch011101010011110110,input1);
	not #50 (output0_branch011101010011110111100,input1);
	not #50 (output0_branch0111010100111101111010,input1);
	and #50 (output0_branch0111010100111101111011100,input0,input0);
	nand #50 (output0_branch011101010011110111101110,output0_branch0111010100111101111011100,input3);
	not #50 (output0_branch01110101001111011110111110100,input1);
	nand #50 (output0_branch0111010100111101111011111010100,input0,input4);
	not #50 (output0_branch01110101001111011110111110101010,input1);
	not #50 (output0_branch011101010011110111101111101010110,input1);
	not #50 (output0_branch0111010100111101111011111010101110,input1);
	not #50 (output0_branch01110101001111011110111110101011110,input1);
	and #50 (output0_branch011101010011110111101111101010111110,input0,input0);
	and #50 (output0_branch01110101001111011110111110101011111100,input0,input0);
	nand #50 (output0_branch0111010100111101111011111010101111110,output0_branch01110101001111011110111110101011111100,input3);
	and #50 (output0_branch0111010100111101111011111010101111111100010000,input0,input0);
	nand #50 (output0_branch011101010011110111101111101010111111110001000,output0_branch0111010100111101111011111010101111111100010000,input3);
	not #50 (output0_branch01110101001111011110111110101011111111000100110100,input1);
	and #50 (output0_branch0111010100111101111011111010101111111100010011010,output0_branch01110101001111011110111110101011111111000100110100,input1);
	not #50 (output0_branch01110101001111011110111110101011111111000100110110100,input1);
	nand #50 (output0_branch0111010100111101111011111010101111111100010011011010100,input0,input4);
	not #50 (output0_branch01110101001111011110111110101011111111000100110110101010,input1);
	not #50 (output0_branch011101010011110111101111101010111111110001001101101010110,input1);
	and #50 (output0_branch011101010011110111101111101010111111110001001101101010111100,input0,input0);
	nand #50 (output0_branch01110101001111011110111110101011111111000100110110101011110,output0_branch011101010011110111101111101010111111110001001101101010111100,input3);
	not #50 (output0_branch0111010100111101111011111010101111111100010011011010101111110100,input1);
	not #50 (output0_branch011101010011110111101111101010111111110001001101101010111111010100,input1);
	xor #50 (output0_branch01110101001111011110111110101011111111000100110110101011111101010,output0_branch011101010011110111101111101010111111110001001101101010111111010100,input3);
	xor #50 (output0_branch0111010100111101111011111010101111111100010011011010101111110101,output0_branch01110101001111011110111110101011111111000100110110101011111101010,input3);
	and #50 (output0_branch011101010011110111101111101010111111110001001101101010111111010,output0_branch0111010100111101111011111010101111111100010011011010101111110100,output0_branch0111010100111101111011111010101111111100010011011010101111110101);
	xor #50 (output0_branch01110101001111011110111110101011111111000100110110101011111101,output0_branch011101010011110111101111101010111111110001001101101010111111010,input0);
	and #50 (output0_branch0111010100111101111011111010101111111100010011011010101111110,input0,output0_branch01110101001111011110111110101011111111000100110110101011111101);
	or #50 (output0_branch011101010011110111101111101010111111110001001101101010111111,output0_branch0111010100111101111011111010101111111100010011011010101111110,input0);
	xor #50 (output0_branch01110101001111011110111110101011111111000100110110101011111,input2,output0_branch011101010011110111101111101010111111110001001101101010111111);
	and #50 (output0_branch0111010100111101111011111010101111111100010011011010101111,output0_branch01110101001111011110111110101011111111000100110110101011110,output0_branch01110101001111011110111110101011111111000100110110101011111);
	or #50 (output0_branch011101010011110111101111101010111111110001001101101010111,input0,output0_branch0111010100111101111011111010101111111100010011011010101111);
	and #50 (output0_branch01110101001111011110111110101011111111000100110110101011,output0_branch011101010011110111101111101010111111110001001101101010110,output0_branch011101010011110111101111101010111111110001001101101010111);
	and #50 (output0_branch0111010100111101111011111010101111111100010011011010101,output0_branch01110101001111011110111110101011111111000100110110101010,output0_branch01110101001111011110111110101011111111000100110110101011);
	xor #50 (output0_branch011101010011110111101111101010111111110001001101101010,output0_branch0111010100111101111011111010101111111100010011011010100,output0_branch0111010100111101111011111010101111111100010011011010101);
	xor #50 (output0_branch01110101001111011110111110101011111111000100110110101,output0_branch011101010011110111101111101010111111110001001101101010,input3);
	and #50 (output0_branch0111010100111101111011111010101111111100010011011010,output0_branch01110101001111011110111110101011111111000100110110100,output0_branch01110101001111011110111110101011111111000100110110101);
	xor #50 (output0_branch011101010011110111101111101010111111110001001101101,output0_branch0111010100111101111011111010101111111100010011011010,input0);
	and #50 (output0_branch01110101001111011110111110101011111111000100110110,input0,output0_branch011101010011110111101111101010111111110001001101101);
	or #50 (output0_branch0111010100111101111011111010101111111100010011011,output0_branch01110101001111011110111110101011111111000100110110,input0);
	xor #50 (output0_branch011101010011110111101111101010111111110001001101,output0_branch0111010100111101111011111010101111111100010011010,output0_branch0111010100111101111011111010101111111100010011011);
	and #50 (output0_branch01110101001111011110111110101011111111000100110,input0,output0_branch011101010011110111101111101010111111110001001101);
	or #50 (output0_branch0111010100111101111011111010101111111100010011,output0_branch01110101001111011110111110101011111111000100110,input0);
	xor #50 (output0_branch011101010011110111101111101010111111110001001,input2,output0_branch0111010100111101111011111010101111111100010011);
	and #50 (output0_branch01110101001111011110111110101011111111000100,output0_branch011101010011110111101111101010111111110001000,output0_branch011101010011110111101111101010111111110001001);
	nand #50 (output0_branch0111010100111101111011111010101111111100010100,input0,input4);
	not #50 (output0_branch01110101001111011110111110101011111111000101010,input1);
	not #50 (output0_branch011101010011110111101111101010111111110001010110,input1);
	or #50 (output0_branch011101010011110111101111101010111111110001010111,input0,input0);
	and #50 (output0_branch01110101001111011110111110101011111111000101011,output0_branch011101010011110111101111101010111111110001010110,output0_branch011101010011110111101111101010111111110001010111);
	and #50 (output0_branch0111010100111101111011111010101111111100010101,output0_branch01110101001111011110111110101011111111000101010,output0_branch01110101001111011110111110101011111111000101011);
	xor #50 (output0_branch011101010011110111101111101010111111110001010,output0_branch0111010100111101111011111010101111111100010100,output0_branch0111010100111101111011111010101111111100010101);
	xor #50 (output0_branch01110101001111011110111110101011111111000101,output0_branch011101010011110111101111101010111111110001010,input3);
	and #50 (output0_branch0111010100111101111011111010101111111100010,output0_branch01110101001111011110111110101011111111000100,output0_branch01110101001111011110111110101011111111000101);
	xor #50 (output0_branch011101010011110111101111101010111111110001,output0_branch0111010100111101111011111010101111111100010,input0);
	and #50 (output0_branch01110101001111011110111110101011111111000,input0,output0_branch011101010011110111101111101010111111110001);
	or #50 (output0_branch0111010100111101111011111010101111111100,output0_branch01110101001111011110111110101011111111000,input0);
	and #50 (output0_branch01110101001111011110111110101011111111010000,input0,input0);
	nand #50 (output0_branch0111010100111101111011111010101111111101000,output0_branch01110101001111011110111110101011111111010000,input3);
	not #50 (output0_branch011101010011110111101111101010111111110100110100,input1);
	and #50 (output0_branch01110101001111011110111110101011111111010011010,output0_branch011101010011110111101111101010111111110100110100,input1);
	not #50 (output0_branch011101010011110111101111101010111111110100110110100,input1);
	nand #50 (output0_branch01110101001111011110111110101011111111010011011010100,input0,input4);
	not #50 (output0_branch011101010011110111101111101010111111110100110110101010,input1);
	not #50 (output0_branch0111010100111101111011111010101111111101001101101010110,input1);
	and #50 (output0_branch0111010100111101111011111010101111111101001101101010111100,input0,input0);
	nand #50 (output0_branch011101010011110111101111101010111111110100110110101011110,output0_branch0111010100111101111011111010101111111101001101101010111100,input3);
	not #50 (output0_branch01110101001111011110111110101011111111010011011010101111110100,input1);
	xor #50 (output0_branch01110101001111011110111110101011111111010011011010101111110101,input1,input3);
	and #50 (output0_branch0111010100111101111011111010101111111101001101101010111111010,output0_branch01110101001111011110111110101011111111010011011010101111110100,output0_branch01110101001111011110111110101011111111010011011010101111110101);
	xor #50 (output0_branch011101010011110111101111101010111111110100110110101011111101,output0_branch0111010100111101111011111010101111111101001101101010111111010,input0);
	and #50 (output0_branch01110101001111011110111110101011111111010011011010101111110,input0,output0_branch011101010011110111101111101010111111110100110110101011111101);
	or #50 (output0_branch0111010100111101111011111010101111111101001101101010111111,output0_branch01110101001111011110111110101011111111010011011010101111110,input0);
	xor #50 (output0_branch011101010011110111101111101010111111110100110110101011111,input2,output0_branch0111010100111101111011111010101111111101001101101010111111);
	and #50 (output0_branch01110101001111011110111110101011111111010011011010101111,output0_branch011101010011110111101111101010111111110100110110101011110,output0_branch011101010011110111101111101010111111110100110110101011111);
	or #50 (output0_branch0111010100111101111011111010101111111101001101101010111,input0,output0_branch01110101001111011110111110101011111111010011011010101111);
	and #50 (output0_branch011101010011110111101111101010111111110100110110101011,output0_branch0111010100111101111011111010101111111101001101101010110,output0_branch0111010100111101111011111010101111111101001101101010111);
	and #50 (output0_branch01110101001111011110111110101011111111010011011010101,output0_branch011101010011110111101111101010111111110100110110101010,output0_branch011101010011110111101111101010111111110100110110101011);
	xor #50 (output0_branch0111010100111101111011111010101111111101001101101010,output0_branch01110101001111011110111110101011111111010011011010100,output0_branch01110101001111011110111110101011111111010011011010101);
	xor #50 (output0_branch011101010011110111101111101010111111110100110110101,output0_branch0111010100111101111011111010101111111101001101101010,input3);
	and #50 (output0_branch01110101001111011110111110101011111111010011011010,output0_branch011101010011110111101111101010111111110100110110100,output0_branch011101010011110111101111101010111111110100110110101);
	xor #50 (output0_branch0111010100111101111011111010101111111101001101101,output0_branch01110101001111011110111110101011111111010011011010,input0);
	and #50 (output0_branch011101010011110111101111101010111111110100110110,input0,output0_branch0111010100111101111011111010101111111101001101101);
	or #50 (output0_branch01110101001111011110111110101011111111010011011,output0_branch011101010011110111101111101010111111110100110110,input0);
	xor #50 (output0_branch0111010100111101111011111010101111111101001101,output0_branch01110101001111011110111110101011111111010011010,output0_branch01110101001111011110111110101011111111010011011);
	and #50 (output0_branch011101010011110111101111101010111111110100110,input0,output0_branch0111010100111101111011111010101111111101001101);
	or #50 (output0_branch01110101001111011110111110101011111111010011,output0_branch011101010011110111101111101010111111110100110,input0);
	xor #50 (output0_branch0111010100111101111011111010101111111101001,input2,output0_branch01110101001111011110111110101011111111010011);
	and #50 (output0_branch011101010011110111101111101010111111110100,output0_branch0111010100111101111011111010101111111101000,output0_branch0111010100111101111011111010101111111101001);
	nand #50 (output0_branch01110101001111011110111110101011111111010100,input0,input4);
	not #50 (output0_branch011101010011110111101111101010111111110101010,input1);
	not #50 (output0_branch0111010100111101111011111010101111111101010110,input1);
	or #50 (output0_branch0111010100111101111011111010101111111101010111,input0,input0);
	and #50 (output0_branch011101010011110111101111101010111111110101011,output0_branch0111010100111101111011111010101111111101010110,output0_branch0111010100111101111011111010101111111101010111);
	and #50 (output0_branch01110101001111011110111110101011111111010101,output0_branch011101010011110111101111101010111111110101010,output0_branch011101010011110111101111101010111111110101011);
	xor #50 (output0_branch0111010100111101111011111010101111111101010,output0_branch01110101001111011110111110101011111111010100,output0_branch01110101001111011110111110101011111111010101);
	xor #50 (output0_branch011101010011110111101111101010111111110101,output0_branch0111010100111101111011111010101111111101010,input3);
	and #50 (output0_branch01110101001111011110111110101011111111010,output0_branch011101010011110111101111101010111111110100,output0_branch011101010011110111101111101010111111110101);
	xor #50 (output0_branch0111010100111101111011111010101111111101,output0_branch01110101001111011110111110101011111111010,input0);
	and #50 (output0_branch011101010011110111101111101010111111110,output0_branch0111010100111101111011111010101111111100,output0_branch0111010100111101111011111010101111111101);
	or #50 (output0_branch01110101001111011110111110101011111111,output0_branch011101010011110111101111101010111111110,input0);
	xor #50 (output0_branch0111010100111101111011111010101111111,input2,output0_branch01110101001111011110111110101011111111);
	and #50 (output0_branch011101010011110111101111101010111111,output0_branch0111010100111101111011111010101111110,output0_branch0111010100111101111011111010101111111);
	or #50 (output0_branch01110101001111011110111110101011111,output0_branch011101010011110111101111101010111110,output0_branch011101010011110111101111101010111111);
	and #50 (output0_branch0111010100111101111011111010101111,output0_branch01110101001111011110111110101011110,output0_branch01110101001111011110111110101011111);
	and #50 (output0_branch011101010011110111101111101010111,output0_branch0111010100111101111011111010101110,output0_branch0111010100111101111011111010101111);
	and #50 (output0_branch01110101001111011110111110101011,output0_branch011101010011110111101111101010110,output0_branch011101010011110111101111101010111);
	and #50 (output0_branch0111010100111101111011111010101,output0_branch01110101001111011110111110101010,output0_branch01110101001111011110111110101011);
	xor #50 (output0_branch011101010011110111101111101010,output0_branch0111010100111101111011111010100,output0_branch0111010100111101111011111010101);
	xor #50 (output0_branch01110101001111011110111110101,output0_branch011101010011110111101111101010,input3);
	and #50 (output0_branch0111010100111101111011111010,output0_branch01110101001111011110111110100,output0_branch01110101001111011110111110101);
	xor #50 (output0_branch011101010011110111101111101,output0_branch0111010100111101111011111010,input0);
	and #50 (output0_branch01110101001111011110111110,input0,output0_branch011101010011110111101111101);
	or #50 (output0_branch0111010100111101111011111,output0_branch01110101001111011110111110,input0);
	xor #50 (output0_branch011101010011110111101111,input2,output0_branch0111010100111101111011111);
	and #50 (output0_branch01110101001111011110111,output0_branch011101010011110111101110,output0_branch011101010011110111101111);
	or #50 (output0_branch0111010100111101111011,input0,output0_branch01110101001111011110111);
	and #50 (output0_branch011101010011110111101,output0_branch0111010100111101111010,output0_branch0111010100111101111011);
	and #50 (output0_branch01110101001111011110,output0_branch011101010011110111100,output0_branch011101010011110111101);
	and #50 (output0_branch0111010100111101111,output0_branch01110101001111011110,input3);
	or #50 (output0_branch011101010011110111,input0,output0_branch0111010100111101111);
	and #50 (output0_branch01110101001111011,output0_branch011101010011110110,output0_branch011101010011110111);
	and #50 (output0_branch0111010100111101,output0_branch01110101001111010,output0_branch01110101001111011);
	xor #50 (output0_branch011101010011110,input3,output0_branch0111010100111101);
	and #50 (output0_branch01110101001111,output0_branch011101010011110,input3);
	or #50 (output0_branch0111010100111,input0,output0_branch01110101001111);
	and #50 (output0_branch011101010011,output0_branch0111010100110,output0_branch0111010100111);
	and #50 (output0_branch01110101001,output0_branch011101010010,output0_branch011101010011);
	xor #50 (output0_branch0111010100,output0_branch01110101000,output0_branch01110101001);
	not #50 (output0_branch01110101010,input1);
	not #50 (output0_branch011101010110,input1);
	not #50 (output0_branch01110101011110010100,input1);
	not #50 (output0_branch011101010111100101010000,input1);
	not #50 (output0_branch0111010101111001010100010,input1);
	not #50 (output0_branch011101010111100101010001110010100,input1);
	nand #50 (output0_branch01110101011110010101000111001010100,input0,input4);
	not #50 (output0_branch011101010111100101010001110010101010,input1);
	not #50 (output0_branch0111010101111001010100011100101010110,input1);
	and #50 (output0_branch0111010101111001010100011100101010111100,input0,input0);
	nand #50 (output0_branch011101010111100101010001110010101011110,output0_branch0111010101111001010100011100101010111100,input3);
	not #50 (output0_branch0111010101111001010100011100101010111111010000,input1);
	nand #50 (output0_branch011101010111100101010001110010101011111101000100,input0,input4);
	not #50 (output0_branch0111010101111001010100011100101010111111010001010,input1);
	not #50 (output0_branch01110101011110010101000111001010101111110100010110,input1);
	and #50 (output0_branch01110101011110010101000111001010101111110100010111100,input0,input0);
	nand #50 (output0_branch0111010101111001010100011100101010111111010001011110,output0_branch01110101011110010101000111001010101111110100010111100,input3);
	or #50 (output0_branch01110101011110010101000111001010101111110100010111111010,input1,input1);
	and #50 (output0_branch0111010101111001010100011100101010111111010001011111101,output0_branch01110101011110010101000111001010101111110100010111111010,input2);
	and #50 (output0_branch011101010111100101010001110010101011111101000101111110,input0,output0_branch0111010101111001010100011100101010111111010001011111101);
	or #50 (output0_branch01110101011110010101000111001010101111110100010111111,output0_branch011101010111100101010001110010101011111101000101111110,input0);
	xor #50 (output0_branch0111010101111001010100011100101010111111010001011111,input2,output0_branch01110101011110010101000111001010101111110100010111111);
	and #50 (output0_branch011101010111100101010001110010101011111101000101111,output0_branch0111010101111001010100011100101010111111010001011110,output0_branch0111010101111001010100011100101010111111010001011111);
	or #50 (output0_branch01110101011110010101000111001010101111110100010111,input0,output0_branch011101010111100101010001110010101011111101000101111);
	and #50 (output0_branch0111010101111001010100011100101010111111010001011,output0_branch01110101011110010101000111001010101111110100010110,output0_branch01110101011110010101000111001010101111110100010111);
	and #50 (output0_branch011101010111100101010001110010101011111101000101,output0_branch0111010101111001010100011100101010111111010001010,output0_branch0111010101111001010100011100101010111111010001011);
	xor #50 (output0_branch01110101011110010101000111001010101111110100010,output0_branch011101010111100101010001110010101011111101000100,output0_branch011101010111100101010001110010101011111101000101);
	xor #50 (output0_branch0111010101111001010100011100101010111111010001,output0_branch01110101011110010101000111001010101111110100010,input3);
	and #50 (output0_branch011101010111100101010001110010101011111101000,output0_branch0111010101111001010100011100101010111111010000,output0_branch0111010101111001010100011100101010111111010001);
	xor #50 (output0_branch01110101011110010101000111001010101111110100,output0_branch011101010111100101010001110010101011111101000,input0);
	nand #50 (output0_branch0111010101111001010100011100101010111111010100,input0,input4);
	not #50 (output0_branch01110101011110010101000111001010101111110101010,input1);
	not #50 (output0_branch0111010101111001010100011100101010111111010101100,input4);
	not #50 (output0_branch011101010111100101010001110010101011111101010110,output0_branch0111010101111001010100011100101010111111010101100);
	or #50 (output0_branch011101010111100101010001110010101011111101010111,input0,input4);
	and #50 (output0_branch01110101011110010101000111001010101111110101011,output0_branch011101010111100101010001110010101011111101010110,output0_branch011101010111100101010001110010101011111101010111);
	and #50 (output0_branch0111010101111001010100011100101010111111010101,output0_branch01110101011110010101000111001010101111110101010,output0_branch01110101011110010101000111001010101111110101011);
	xor #50 (output0_branch011101010111100101010001110010101011111101010,output0_branch0111010101111001010100011100101010111111010100,output0_branch0111010101111001010100011100101010111111010101);
	xor #50 (output0_branch01110101011110010101000111001010101111110101,output0_branch011101010111100101010001110010101011111101010,input3);
	and #50 (output0_branch0111010101111001010100011100101010111111010,output0_branch01110101011110010101000111001010101111110100,output0_branch01110101011110010101000111001010101111110101);
	xor #50 (output0_branch011101010111100101010001110010101011111101,output0_branch0111010101111001010100011100101010111111010,input0);
	and #50 (output0_branch01110101011110010101000111001010101111110,input0,output0_branch011101010111100101010001110010101011111101);
	or #50 (output0_branch0111010101111001010100011100101010111111,output0_branch01110101011110010101000111001010101111110,input0);
	xor #50 (output0_branch011101010111100101010001110010101011111,input2,output0_branch0111010101111001010100011100101010111111);
	and #50 (output0_branch01110101011110010101000111001010101111,output0_branch011101010111100101010001110010101011110,output0_branch011101010111100101010001110010101011111);
	or #50 (output0_branch0111010101111001010100011100101010111,input0,output0_branch01110101011110010101000111001010101111);
	and #50 (output0_branch011101010111100101010001110010101011,output0_branch0111010101111001010100011100101010110,output0_branch0111010101111001010100011100101010111);
	and #50 (output0_branch01110101011110010101000111001010101,output0_branch011101010111100101010001110010101010,output0_branch011101010111100101010001110010101011);
	xor #50 (output0_branch0111010101111001010100011100101010,output0_branch01110101011110010101000111001010100,output0_branch01110101011110010101000111001010101);
	xor #50 (output0_branch011101010111100101010001110010101,output0_branch0111010101111001010100011100101010,input3);
	and #50 (output0_branch01110101011110010101000111001010,output0_branch011101010111100101010001110010100,output0_branch011101010111100101010001110010101);
	xor #50 (output0_branch0111010101111001010100011100101,output0_branch01110101011110010101000111001010,input0);
	and #50 (output0_branch011101010111100101010001110010,input0,output0_branch0111010101111001010100011100101);
	or #50 (output0_branch01110101011110010101000111001,output0_branch011101010111100101010001110010,input0);
	xor #50 (output0_branch0111010101111001010100011100,input2,output0_branch01110101011110010101000111001);
	not #50 (output0_branch011101010111100101010001110,output0_branch0111010101111001010100011100);
	not #50 (output0_branch0111010101111001010100011110,input1);
	and #50 (output0_branch01110101011110010101000111110100,input0,input0);
	nand #50 (output0_branch0111010101111001010100011111010,output0_branch01110101011110010101000111110100,input3);
	and #50 (output0_branch011101010111100101010001111101,output0_branch0111010101111001010100011111010,input3);
	or #50 (output0_branch01110101011110010101000111110,input0,output0_branch011101010111100101010001111101);
	and #50 (output0_branch0111010101111001010100011111100,input0,input0);
	nand #50 (output0_branch011101010111100101010001111110,output0_branch0111010101111001010100011111100,input3);
	and #50 (output0_branch01110101011110010101000111111,output0_branch011101010111100101010001111110,input3);
	or #50 (output0_branch0111010101111001010100011111,output0_branch01110101011110010101000111110,output0_branch01110101011110010101000111111);
	and #50 (output0_branch011101010111100101010001111,output0_branch0111010101111001010100011110,output0_branch0111010101111001010100011111);
	and #50 (output0_branch01110101011110010101000111,output0_branch011101010111100101010001110,output0_branch011101010111100101010001111);
	or #50 (output0_branch0111010101111001010100011,input0,output0_branch01110101011110010101000111);
	and #50 (output0_branch011101010111100101010001,output0_branch0111010101111001010100010,output0_branch0111010101111001010100011);
	and #50 (output0_branch01110101011110010101000,output0_branch011101010111100101010000,output0_branch011101010111100101010001);
	nand #50 (output0_branch0111010101111001010100,output0_branch01110101011110010101000,input4);
	not #50 (output0_branch011101010111100101010110,input1);
	and #50 (output0_branch011101010111100101010111100,input0,input0);
	nand #50 (output0_branch01110101011110010101011110,output0_branch011101010111100101010111100,input3);
	and #50 (output0_branch0111010101111001010101111,output0_branch01110101011110010101011110,input3);
	or #50 (output0_branch011101010111100101010111,input0,output0_branch0111010101111001010101111);
	and #50 (output0_branch01110101011110010101011,output0_branch011101010111100101010110,output0_branch011101010111100101010111);
	and #50 (output0_branch0111010101111001010101,input0,output0_branch01110101011110010101011);
	xor #50 (output0_branch011101010111100101010,output0_branch0111010101111001010100,output0_branch0111010101111001010101);
	xor #50 (output0_branch01110101011110010101,output0_branch011101010111100101010,input3);
	and #50 (output0_branch0111010101111001010,output0_branch01110101011110010100,output0_branch01110101011110010101);
	xor #50 (output0_branch011101010111100101,output0_branch0111010101111001010,input0);
	and #50 (output0_branch01110101011110010,input0,output0_branch011101010111100101);
	or #50 (output0_branch0111010101111001,output0_branch01110101011110010,input0);
	xor #50 (output0_branch011101010111100,input2,output0_branch0111010101111001);
	nand #50 (output0_branch01110101011110,output0_branch011101010111100,input3);
	and #50 (output0_branch0111010101111,output0_branch01110101011110,input3);
	or #50 (output0_branch011101010111,input0,output0_branch0111010101111);
	and #50 (output0_branch01110101011,output0_branch011101010110,output0_branch011101010111);
	and #50 (output0_branch0111010101,output0_branch01110101010,output0_branch01110101011);
	xor #50 (output0_branch011101010,output0_branch0111010100,output0_branch0111010101);
	xor #50 (output0_branch01110101,output0_branch011101010,input0);
	and #50 (output0_branch0111010,output0_branch01110100,output0_branch01110101);
	xor #50 (output0_branch011101,output0_branch0111010,input0);
	and #50 (output0_branch01110,input0,output0_branch011101);
	or #50 (output0_branch0111,output0_branch01110,input0);
	xor #50 (output0_branch011,input2,output0_branch0111);
	and #50 (output0_branch01,output0_branch010,output0_branch011);
	or #50 (output0,input0,output0_branch01);

	and #50 (output1_branch01000,input0,input2);
	nand #50 (output1_branch01001,input1,input1);
	xor #50 (output1_branch0100,output1_branch01000,output1_branch01001);
	not #50 (output1_branch010,output1_branch0100);
	or #50 (output1_branch01111,input0,input1);
	or #50 (output1_branch0111,input0,output1_branch01111);
	or #50 (output1_branch011,input1,output1_branch0111);
	or #50 (output1_branch01,output1_branch010,output1_branch011);
	or #50 (output1,input0,output1_branch01);

	nand #50 (output2,input0,input0);

	not #50 (output3,input1);


endmodule