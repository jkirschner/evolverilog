module andTest(output0,input0,input1);

	output output0;
	input input0,input1;

	wire output0;

	xor #50 (output0,input0,input0);

endmodule