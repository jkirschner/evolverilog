module andTest(out,A,B);

    output out;
    input A,B;

    and #50 (out,A,B);

endmodule
